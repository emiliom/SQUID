netcdf SQUID_all {
dimensions:
	trajectory = 18 ;
	obs = 234 ;
	z = 2001 ;
	trid_len = 6 ;
variables:
	int trajectory(trajectory) ;
		trajectory:long_name = "Unique identifier for each feature instance" ;
		trajectory:cf_role = "trajectory_id" ;
		trajectory:comment = "ID number of Float-Deployment pair" ;
	double time(obs, trajectory) ;
		time:_FillValue = -9999. ;
		time:long_name = "Time, UTC" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00 0:00" ;
		time:calendar = "Julian" ;
		time:axis = "T" ;
	double lat(obs, trajectory) ;
		lat:_FillValue = -9999. ;
		lat:long_name = "mean latitude of EM-APEX profiles" ;
		lat:standard_name = "latitude" ;
		lat:units = "degree_north" ;
		lat:axis = "Y" ;
		lat:valid_min = "-34.012" ;
		lat:valid_max = "37.1694" ;
		lat:comment = "Mean latitude during each float dive" ;
		lat:Coordinates = "time lat lon" ;
	double lon(obs, trajectory) ;
		lon:_FillValue = -9999. ;
		lon:long_name = "mean longitude of EM-APEX profiles" ;
		lon:standard_name = "longitude" ;
		lon:units = "degree_east" ;
		lon:axis = "X" ;
		lon:valid_min = "-125.105" ;
		lon:valid_max = "93.4306" ;
		lon:comment = "Mean longitude during each float dive" ;
		lon:Coordinates = "time lat lon" ;
	double depth(z, obs, trajectory) ;
		depth:_FillValue = -9999. ;
		depth:long_name = "depths of gridded EM-APEX profiles" ;
		depth:standard_name = "depth" ;
		depth:units = "meters [m]" ;
		depth:axis = "Z" ;
		depth:positive = "down" ;
		depth:valid_min = "0" ;
		depth:valid_max = "-2000" ;
		depth:comment = "Profile depths interpolated to common grid" ;
	double T(z, obs, trajectory) ;
		T:_FillValue = -9999. ;
		T:long_name = "gridded EM-APEX temperature" ;
		T:standard_name = "sea_water_temperature" ;
		T:units = "Kelvin" ;
		T:coordinates = "time lat lon z" ;
		T:platform_variable = "EM_APEX" ;
		T:instrument = "thermistor" ;
	double S(z, obs, trajectory) ;
		S:_FillValue = -9999. ;
		S:long_name = "gridded EM-APEX salinity" ;
		S:standard_name = "sea_water_salinity" ;
		S:units = "1e-3" ;
		S:coordinates = "time lat lon z" ;
		S:platform_variable = "EM_APEX" ;
		S:comment = "Units are standard psu. The units refered to in Units attribute refer to the CF Convention for standard name and units." ;
	double P(z, obs, trajectory) ;
		P:_FillValue = -9999. ;
		P:long_name = "gridded EM-APEX pressure derived from depth and latitude" ;
		P:standard_name = "sea_water_pressure" ;
		P:units = "decibar" ;
		P:coordinates = "time lat lon z" ;
		P:platform_variable = "EM_APEX" ;
	double U(z, obs, trajectory) ;
		U:_FillValue = -9999. ;
		U:long_name = "gridded EM-APEX east velocity component" ;
		U:standard_name = "eastward_sea_water_velocity" ;
		U:units = "meter per second" ;
		U:coordinates = "time lat lon z" ;
		U:platform_variable = "EM_APEX" ;
		U:instrument = "EM-APEX" ;
	double V(z, obs, trajectory) ;
		V:_FillValue = -9999. ;
		V:long_name = "gridded EM-APEX north velocity component" ;
		V:standard_name = "northward_sea_water_velocity" ;
		V:units = "meter per second" ;
		V:coordinates = "time lat lon z" ;
		V:platform_variable = "EM_APEX" ;
		V:instrument = "EM-APEX" ;
	double chi1(z, obs, trajectory) ;
		chi1:_FillValue = -9999. ;
		chi1:long_name = "temperature_variance_dissipation" ;
		chi1:units = "degree Celsius square per second" ;
		chi1:coordinates = "time lat lon z" ;
		chi1:platform_variable = "EM_APEX" ;
		chi1:comment = "Rate of dissipation of temperature variance measured by Probe 1" ;
	double chi2(z, obs, trajectory) ;
		chi2:_FillValue = -9999. ;
		chi2:long_name = "temperature_variance_dissipation" ;
		chi2:units = "degree Celsius square per second" ;
		chi2:coordinates = "time lat lon z" ;
		chi2:platform_variable = "EM_APEX" ;
		chi2:comment = "Rate of dissipation of temperature variance measured by Probe 2" ;
	double ptime(z, obs, trajectory) ;
		ptime:_FillValue = -9999. ;
		ptime:long_name = "time_along_profile" ;
		ptime:units = "seconds since 1970-01-01 00:00:00 0:00" ;
		ptime:calendar = "Julian" ;
		ptime:coordinates = "time lat lon z" ;
		ptime:platform_variable = "EM_APEX" ;
	double U0(obs, trajectory) ;
		U0:_FillValue = -9999. ;
		U0:long_name = "Drift eastward velocity of a float while at surface" ;
		U0:standard_name = "surface eastward velocity" ;
		U0:units = "meter per second" ;
		U0:Coordinates = "time lat lon" ;
	double V0(obs, trajectory) ;
		V0:_FillValue = -9999. ;
		V0:long_name = "Drift northward velocity of a float while at surface" ;
		V0:standard_name = "surface northward velocity" ;
		V0:units = "meter per second" ;
		V0:Coordinates = "time lat lon" ;
	int flid(trajectory) ;
		flid:long_name = "EM-APEX float id number" ;
		flid:standard_name = "Float id number" ;
	char trid(trid_len, trajectory) ;
		trid:long_name = "Trajectory id" ;
		trid:comment = "A 2-dimensional character array representing a unique trajectory id string per float deployment. The rendering of this trajectory id is dependent on the software used to read the netcdfs. If the trajectory id does not look like a composition of a float number and characters (e.g. \'f9436\', \'7805s2\'), try to compose the trajectory id string by concatenating the characters over the trid_len dimension" ;
	int pid(obs, trajectory) ;
		pid:_FillValue = -9999 ;
		pid:long_name = "Profile id number" ;
		pid:comment = "Profile number, where a profile consist of a full down + up cycle" ;
	int hpid(obs, trajectory) ;
		hpid:_FillValue = -9999 ;
		hpid:long_name = "Half-profile id number" ;
		hpid:comment = "A Half profile consist of either a down or up profile. Odd number are down-profiles, even numbers are up-profiles" ;
	int depl(trajectory) ;
		depl:long_name = "Deployment number of a float" ;
		depl:standard_name = "deployment" ;
		depl:comment = "Deployment number within an experiment. An experiment can have a single deployment or multiple deployments where all or part of the float array are deployed. " ;
	double EM-APEX ;
		EM-APEX:_FillValue = -9999. ;
		EM-APEX:long_name = "EM-APEX" ;
		EM-APEX:wmo_code = "" ;

// global attributes:
		:ncei_template_version = "NCEI_NetCDF_TrajectoryProfile_Incomplete_Template_v2.0" ;
		:featureType = "trajectoryProfile" ;
		:title = "T, S, U, V and derived quantities measured by EM-APEX during SQUIDexperiment" ;
		:summary = "T, S, potential density, N^2, U, V, u_z, and v_z measured by EM-APEX float and interpolated onto a common depth grid" ;
		:Conventions = "CF-1.6, ACDD-1.3" ;
		:acknowledgments = "NOPP Global Internal Wave Project. Funding from the National Science Foundation (OCE-2232796)" ;
		:date_created = "19-Mar-2024 04:49:52" ;
		:creator_name = "James Girton, Aurelie Moulin" ;
		:creator_email = "girton@uw.edu, amoulin@uw.edu" ;
		:Institution = "Applied Physics Laboratory - University of Washington" ;
		:geospatial_lat_min = "-59.1682 (>0, N; <0, S)" ;
		:geospatial_lat_max = "40.8682 (>0, N; <0, S)" ;
		:geospatial_lon_min = "-127.4163 (>0, E; <0, W)" ;
		:geospatial_lon_max = "155.869 (>0, E; <0, W)" ;
		:vertical_min = -2000. ;
		:vertical_max = -0. ;
		:vertical_positive = "up" ;
		:time_coverage_start = "18-Feb-2023 21:11:05" ;
		:time_coverage_end = "14-Mar-2024 10:19:33" ;
		:sea_name = "Multiple" ;
		:geospatial_lat_units = "degree_north" ;
		:geospatial_lon_units = "degree_east" ;
		:geospatial_vertical_units = "meters" ;
		:platform = "EM-APEX" ;
		:references = "" ;
		:comment = "Deployed from multiple cruises of opportunity worlwide for the Sampling Quantitative Internal Waves Dissipation project (SQUID)starting in Feb 2023. PI: James Girton (girton@uw.edu)" ;
}
